// Raster_Laser_Projector_Video_In.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module Raster_Laser_Projector_Video_In (
		input  wire        clk_clk,                  //          clk.clk
		input  wire        reset_reset_n,            //        reset.reset_n
		input  wire        video_in_TD_CLK27,        //     video_in.TD_CLK27
		input  wire [7:0]  video_in_TD_DATA,         //             .TD_DATA
		input  wire        video_in_TD_HS,           //             .TD_HS
		input  wire        video_in_TD_VS,           //             .TD_VS
		input  wire        video_in_clk27_reset,     //             .clk27_reset
		output wire        video_in_TD_RESET,        //             .TD_RESET
		output wire        video_in_overflow_flag,   //             .overflow_flag
		output wire [31:0] video_in_dma_address,     // video_in_dma.address
		input  wire        video_in_dma_waitrequest, //             .waitrequest
		output wire        video_in_dma_write,       //             .write
		output wire [7:0]  video_in_dma_writedata    //             .writedata
	);

	wire         video_clipper_0_avalon_clipper_source_valid;           // video_clipper_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire   [7:0] video_clipper_0_avalon_clipper_source_data;            // video_clipper_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_clipper_0_avalon_clipper_source_ready;           // video_scaler_0:stream_in_ready -> video_clipper_0:stream_out_ready
	wire         video_clipper_0_avalon_clipper_source_startofpacket;   // video_clipper_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_clipper_0_avalon_clipper_source_endofpacket;     // video_clipper_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         video_csc_avalon_csc_source_valid;                     // video_csc:stream_out_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] video_csc_avalon_csc_source_data;                      // video_csc:stream_out_data -> video_rgb_resampler_0:stream_in_data
	wire         video_csc_avalon_csc_source_ready;                     // video_rgb_resampler_0:stream_in_ready -> video_csc:stream_out_ready
	wire         video_csc_avalon_csc_source_startofpacket;             // video_csc:stream_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_csc_avalon_csc_source_endofpacket;               // video_csc:stream_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_decoder_0_avalon_decoder_source_valid;           // video_decoder_0:stream_out_valid -> video_chroma_resampler_0:stream_in_valid
	wire  [15:0] video_decoder_0_avalon_decoder_source_data;            // video_decoder_0:stream_out_data -> video_chroma_resampler_0:stream_in_data
	wire         video_decoder_0_avalon_decoder_source_ready;           // video_chroma_resampler_0:stream_in_ready -> video_decoder_0:stream_out_ready
	wire         video_decoder_0_avalon_decoder_source_startofpacket;   // video_decoder_0:stream_out_startofpacket -> video_chroma_resampler_0:stream_in_startofpacket
	wire         video_decoder_0_avalon_decoder_source_endofpacket;     // video_decoder_0:stream_out_endofpacket -> video_chroma_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;         // video_rgb_resampler_0:stream_out_valid -> video_clipper_0:stream_in_valid
	wire   [7:0] video_rgb_resampler_0_avalon_rgb_source_data;          // video_rgb_resampler_0:stream_out_data -> video_clipper_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;         // video_clipper_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket; // video_rgb_resampler_0:stream_out_startofpacket -> video_clipper_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;   // video_rgb_resampler_0:stream_out_endofpacket -> video_clipper_0:stream_in_endofpacket
	wire         video_scaler_0_avalon_scaler_source_valid;             // video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire   [7:0] video_scaler_0_avalon_scaler_source_data;              // video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	wire         video_scaler_0_avalon_scaler_source_ready;             // avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	wire         video_scaler_0_avalon_scaler_source_channel;           // video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         video_scaler_0_avalon_scaler_source_startofpacket;     // video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;       // video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                         // avalon_st_adapter:out_0_valid -> video_dma_controller_0:stream_valid
	wire   [7:0] avalon_st_adapter_out_0_data;                          // avalon_st_adapter:out_0_data -> video_dma_controller_0:stream_data
	wire         avalon_st_adapter_out_0_ready;                         // video_dma_controller_0:stream_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                 // avalon_st_adapter:out_0_startofpacket -> video_dma_controller_0:stream_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                   // avalon_st_adapter:out_0_endofpacket -> video_dma_controller_0:stream_endofpacket
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, video_chroma_resampler_0:reset, video_clipper_0:reset, video_csc:reset, video_decoder_0:reset, video_dma_controller_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]

	Raster_Laser_Projector_Video_In_video_chroma_resampler_0 video_chroma_resampler_0 (
		.clk                      (clk_clk),                                             //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (video_decoder_0_avalon_decoder_source_startofpacket), //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (video_decoder_0_avalon_decoder_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_decoder_0_avalon_decoder_source_valid),         //                     .valid
		.stream_in_ready          (video_decoder_0_avalon_decoder_source_ready),         //                     .ready
		.stream_in_data           (video_decoder_0_avalon_decoder_source_data),          //                     .data
		.stream_out_ready         (),                                                    // avalon_chroma_source.ready
		.stream_out_startofpacket (),                                                    //                     .startofpacket
		.stream_out_endofpacket   (),                                                    //                     .endofpacket
		.stream_out_valid         (),                                                    //                     .valid
		.stream_out_data          ()                                                     //                     .data
	);

	Raster_Laser_Projector_Video_In_video_clipper_0 video_clipper_0 (
		.clk                      (clk_clk),                                               //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //                 reset.reset
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (video_clipper_0_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_0_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (video_clipper_0_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_0_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (video_clipper_0_avalon_clipper_source_valid)            //                      .valid
	);

	Raster_Laser_Projector_Video_In_video_csc video_csc (
		.clk                      (clk_clk),                                   //               clk.clk
		.reset                    (rst_controller_reset_out_reset),            //             reset.reset
		.stream_in_startofpacket  (),                                          //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (),                                          //                  .endofpacket
		.stream_in_valid          (),                                          //                  .valid
		.stream_in_ready          (),                                          //                  .ready
		.stream_in_data           (),                                          //                  .data
		.stream_out_ready         (video_csc_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (video_csc_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_csc_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_csc_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (video_csc_avalon_csc_source_data)           //                  .data
	);

	Raster_Laser_Projector_Video_In_video_decoder_0 video_decoder_0 (
		.clk                      (clk_clk),                                             //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                 reset.reset
		.stream_out_ready         (video_decoder_0_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_decoder_0_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_decoder_0_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_decoder_0_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_decoder_0_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_in_TD_CLK27),                                   //    external_interface.export
		.TD_DATA                  (video_in_TD_DATA),                                    //                      .export
		.TD_HS                    (video_in_TD_HS),                                      //                      .export
		.TD_VS                    (video_in_TD_VS),                                      //                      .export
		.clk27_reset              (video_in_clk27_reset),                                //                      .export
		.TD_RESET                 (video_in_TD_RESET),                                   //                      .export
		.overflow_flag            (video_in_overflow_flag)                               //                      .export
	);

	Raster_Laser_Projector_Video_In_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (clk_clk),                               //                      clk.clk
		.reset                (rst_controller_reset_out_reset),        //                    reset.reset
		.stream_data          (avalon_st_adapter_out_0_data),          //          avalon_dma_sink.data
		.stream_startofpacket (avalon_st_adapter_out_0_startofpacket), //                         .startofpacket
		.stream_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //                         .endofpacket
		.stream_valid         (avalon_st_adapter_out_0_valid),         //                         .valid
		.stream_ready         (avalon_st_adapter_out_0_ready),         //                         .ready
		.slave_address        (),                                      // avalon_dma_control_slave.address
		.slave_byteenable     (),                                      //                         .byteenable
		.slave_read           (),                                      //                         .read
		.slave_write          (),                                      //                         .write
		.slave_writedata      (),                                      //                         .writedata
		.slave_readdata       (),                                      //                         .readdata
		.master_address       (video_in_dma_address),                  //        avalon_dma_master.address
		.master_waitrequest   (video_in_dma_waitrequest),              //                         .waitrequest
		.master_write         (video_in_dma_write),                    //                         .write
		.master_writedata     (video_in_dma_writedata)                 //                         .writedata
	);

	Raster_Laser_Projector_Video_In_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                               //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (video_csc_avalon_csc_source_startofpacket),             //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_csc_avalon_csc_source_endofpacket),               //                  .endofpacket
		.stream_in_valid          (video_csc_avalon_csc_source_valid),                     //                  .valid
		.stream_in_ready          (video_csc_avalon_csc_source_ready),                     //                  .ready
		.stream_in_data           (video_csc_avalon_csc_source_data),                      //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)           //                  .data
	);

	Raster_Laser_Projector_Video_In_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),                                             //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (video_clipper_0_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_0_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_0_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_0_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_0_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data),            //                     .data
		.stream_out_channel       (video_scaler_0_avalon_scaler_source_channel)          //                     .channel
	);

	Raster_Laser_Projector_Video_In_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (1),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                    // in_rst_0.reset
		.in_0_data           (video_scaler_0_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (video_scaler_0_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (video_scaler_0_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (video_scaler_0_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                      //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                     //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                     //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),             //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
