-- Raster_Laser_Projector_Subsystem_0.vhd

-- Generated using ACDS version 16.1 200

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Raster_Laser_Projector_Subsystem_0 is
	port (
		clk_clk               : in std_logic := '0'; --           clk.clk
		hsync_ref_clk         : in std_logic := '0'; --     hsync_ref.clk
		hsync_ref_rst_reset_n : in std_logic := '0'; -- hsync_ref_rst.reset_n
		reset_reset_n         : in std_logic := '0'  --         reset.reset_n
	);
end entity Raster_Laser_Projector_Subsystem_0;

architecture rtl of Raster_Laser_Projector_Subsystem_0 is
begin

end architecture rtl; -- of Raster_Laser_Projector_Subsystem_0
