
module Raster_Laser_Projector (
	clk_50mhz_in_clk,
	pixel_clk_clk,
	reset_reset_n);	

	input		clk_50mhz_in_clk;
	output		pixel_clk_clk;
	input		reset_reset_n;
endmodule
