-- Raster_Laser_Projector.vhd

-- Generated using ACDS version 16.1 200

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Raster_Laser_Projector is
	port (
		clk_50mhz_in_clk                                   : in  std_logic                    := '0';             --                         clk_50mhz_in.clk
		pixel_clk_clk                                      : out std_logic;                                       --                            pixel_clk.clk
		reset_reset_n                                      : in  std_logic                    := '0';             --                                reset.reset_n
		video_in_video_in_external_interface_TD_CLK27      : in  std_logic                    := '0';             -- video_in_video_in_external_interface.TD_CLK27
		video_in_video_in_external_interface_TD_DATA       : in  std_logic_vector(7 downto 0) := (others => '0'); --                                     .TD_DATA
		video_in_video_in_external_interface_TD_HS         : in  std_logic                    := '0';             --                                     .TD_HS
		video_in_video_in_external_interface_TD_VS         : in  std_logic                    := '0';             --                                     .TD_VS
		video_in_video_in_external_interface_clk27_reset   : in  std_logic                    := '0';             --                                     .clk27_reset
		video_in_video_in_external_interface_TD_RESET      : out std_logic;                                       --                                     .TD_RESET
		video_in_video_in_external_interface_overflow_flag : out std_logic                                        --                                     .overflow_flag
	);
end entity Raster_Laser_Projector;

architecture rtl of Raster_Laser_Projector is
	component Raster_Laser_Projector_Clock_Generators is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component Raster_Laser_Projector_Clock_Generators;

	component Raster_Laser_Projector_Framebuffer is
		port (
			address     : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(7 downto 0);                     -- readdata
			writedata   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			address2    : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata2  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			freeze      : in  std_logic                     := 'X';             -- freeze
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component Raster_Laser_Projector_Framebuffer;

	component Raster_Laser_Projector_Video_In is
		port (
			clk_clk                                   : in  std_logic                     := 'X';             -- clk
			reset_reset_n                             : in  std_logic                     := 'X';             -- reset_n
			video_in_dma_address                      : out std_logic_vector(31 downto 0);                    -- address
			video_in_dma_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			video_in_dma_write                        : out std_logic;                                        -- write
			video_in_dma_writedata                    : out std_logic_vector(7 downto 0);                     -- writedata
			video_in_external_interface_TD_CLK27      : in  std_logic                     := 'X';             -- TD_CLK27
			video_in_external_interface_TD_DATA       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- TD_DATA
			video_in_external_interface_TD_HS         : in  std_logic                     := 'X';             -- TD_HS
			video_in_external_interface_TD_VS         : in  std_logic                     := 'X';             -- TD_VS
			video_in_external_interface_clk27_reset   : in  std_logic                     := 'X';             -- clk27_reset
			video_in_external_interface_TD_RESET      : out std_logic;                                        -- TD_RESET
			video_in_external_interface_overflow_flag : out std_logic                                         -- overflow_flag
		);
	end component Raster_Laser_Projector_Video_In;

	component Raster_Laser_Projector_X_Axis_Subsystem is
		port (
			clk_clk             : in std_logic := 'X'; -- clk
			hsync_reset_reset_n : in std_logic := 'X'; -- reset_n
			hsync_target_clk    : in std_logic := 'X'; -- clk
			reset_reset_n       : in std_logic := 'X'  -- reset_n
		);
	end component Raster_Laser_Projector_X_Axis_Subsystem;

	component Raster_Laser_Projector_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			Framebuffer_reset1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Video_In_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			Video_In_video_in_dma_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Video_In_video_in_dma_waitrequest              : out std_logic;                                        -- waitrequest
			Video_In_video_in_dma_write                    : in  std_logic                     := 'X';             -- write
			Video_In_video_in_dma_writedata                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			Framebuffer_s1_address                         : out std_logic_vector(18 downto 0);                    -- address
			Framebuffer_s1_write                           : out std_logic;                                        -- write
			Framebuffer_s1_readdata                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			Framebuffer_s1_writedata                       : out std_logic_vector(7 downto 0);                     -- writedata
			Framebuffer_s1_chipselect                      : out std_logic;                                        -- chipselect
			Framebuffer_s1_clken                           : out std_logic                                         -- clken
		);
	end component Raster_Laser_Projector_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clock_generators_c1_clk                     : std_logic;                     -- Clock_Generators:c1 -> X_Axis_Subsystem:hsync_target_clk
	signal video_in_video_in_dma_waitrequest           : std_logic;                     -- mm_interconnect_0:Video_In_video_in_dma_waitrequest -> Video_In:video_in_dma_waitrequest
	signal video_in_video_in_dma_address               : std_logic_vector(31 downto 0); -- Video_In:video_in_dma_address -> mm_interconnect_0:Video_In_video_in_dma_address
	signal video_in_video_in_dma_write                 : std_logic;                     -- Video_In:video_in_dma_write -> mm_interconnect_0:Video_In_video_in_dma_write
	signal video_in_video_in_dma_writedata             : std_logic_vector(7 downto 0);  -- Video_In:video_in_dma_writedata -> mm_interconnect_0:Video_In_video_in_dma_writedata
	signal mm_interconnect_0_framebuffer_s1_chipselect : std_logic;                     -- mm_interconnect_0:Framebuffer_s1_chipselect -> Framebuffer:chipselect
	signal mm_interconnect_0_framebuffer_s1_readdata   : std_logic_vector(7 downto 0);  -- Framebuffer:readdata -> mm_interconnect_0:Framebuffer_s1_readdata
	signal mm_interconnect_0_framebuffer_s1_address    : std_logic_vector(18 downto 0); -- mm_interconnect_0:Framebuffer_s1_address -> Framebuffer:address
	signal mm_interconnect_0_framebuffer_s1_write      : std_logic;                     -- mm_interconnect_0:Framebuffer_s1_write -> Framebuffer:write
	signal mm_interconnect_0_framebuffer_s1_writedata  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Framebuffer_s1_writedata -> Framebuffer:writedata
	signal mm_interconnect_0_framebuffer_s1_clken      : std_logic;                     -- mm_interconnect_0:Framebuffer_s1_clken -> Framebuffer:clken
	signal rst_controller_reset_out_reset              : std_logic;                     -- rst_controller:reset_out -> [Clock_Generators:reset, Framebuffer:reset, mm_interconnect_0:Framebuffer_reset1_reset_bridge_in_reset_reset, mm_interconnect_0:Video_In_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	clock_generators : component Raster_Laser_Projector_Clock_Generators
		port map (
			clk                => clk_50mhz_in_clk,               --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                           --             pll_slave.read
			write              => open,                           --                      .write
			address            => open,                           --                      .address
			readdata           => open,                           --                      .readdata
			writedata          => open,                           --                      .writedata
			c0                 => open,                           --                    c0.clk
			c1                 => clock_generators_c1_clk,        --                    c1.clk
			c2                 => pixel_clk_clk,                  --                    c2.clk
			areset             => open,                           --        areset_conduit.export
			locked             => open,                           --        locked_conduit.export
			scandone           => open,                           --           (terminated)
			scandataout        => open,                           --           (terminated)
			phasedone          => open,                           --           (terminated)
			phasecounterselect => "0000",                         --           (terminated)
			phaseupdown        => '0',                            --           (terminated)
			phasestep          => '0',                            --           (terminated)
			scanclk            => '0',                            --           (terminated)
			scanclkena         => '0',                            --           (terminated)
			scandata           => '0',                            --           (terminated)
			configupdate       => '0'                             --           (terminated)
		);

	framebuffer : component Raster_Laser_Projector_Framebuffer
		port map (
			address     => mm_interconnect_0_framebuffer_s1_address,    --     s1.address
			clken       => mm_interconnect_0_framebuffer_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_framebuffer_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_framebuffer_s1_write,      --       .write
			readdata    => mm_interconnect_0_framebuffer_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_framebuffer_s1_writedata,  --       .writedata
			address2    => open,                                        --     s2.address
			chipselect2 => open,                                        --       .chipselect
			clken2      => open,                                        --       .clken
			write2      => open,                                        --       .write
			readdata2   => open,                                        --       .readdata
			writedata2  => open,                                        --       .writedata
			clk         => clk_50mhz_in_clk,                            --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			freeze      => '0',                                         -- (terminated)
			reset_req   => '0'                                          -- (terminated)
		);

	video_in : component Raster_Laser_Projector_Video_In
		port map (
			clk_clk                                   => clk_50mhz_in_clk,                                   --                         clk.clk
			reset_reset_n                             => reset_reset_n,                                      --                       reset.reset_n
			video_in_dma_address                      => video_in_video_in_dma_address,                      --                video_in_dma.address
			video_in_dma_waitrequest                  => video_in_video_in_dma_waitrequest,                  --                            .waitrequest
			video_in_dma_write                        => video_in_video_in_dma_write,                        --                            .write
			video_in_dma_writedata                    => video_in_video_in_dma_writedata,                    --                            .writedata
			video_in_external_interface_TD_CLK27      => video_in_video_in_external_interface_TD_CLK27,      -- video_in_external_interface.TD_CLK27
			video_in_external_interface_TD_DATA       => video_in_video_in_external_interface_TD_DATA,       --                            .TD_DATA
			video_in_external_interface_TD_HS         => video_in_video_in_external_interface_TD_HS,         --                            .TD_HS
			video_in_external_interface_TD_VS         => video_in_video_in_external_interface_TD_VS,         --                            .TD_VS
			video_in_external_interface_clk27_reset   => video_in_video_in_external_interface_clk27_reset,   --                            .clk27_reset
			video_in_external_interface_TD_RESET      => video_in_video_in_external_interface_TD_RESET,      --                            .TD_RESET
			video_in_external_interface_overflow_flag => video_in_video_in_external_interface_overflow_flag  --                            .overflow_flag
		);

	x_axis_subsystem : component Raster_Laser_Projector_X_Axis_Subsystem
		port map (
			clk_clk             => clk_50mhz_in_clk,        --          clk.clk
			hsync_reset_reset_n => reset_reset_n,           --  hsync_reset.reset_n
			hsync_target_clk    => clock_generators_c1_clk, -- hsync_target.clk
			reset_reset_n       => reset_reset_n            --        reset.reset_n
		);

	mm_interconnect_0 : component Raster_Laser_Projector_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_50mhz_in_clk,                            --                                clk_0_clk.clk
			Framebuffer_reset1_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,              -- Framebuffer_reset1_reset_bridge_in_reset.reset
			Video_In_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,              --     Video_In_reset_reset_bridge_in_reset.reset
			Video_In_video_in_dma_address                  => video_in_video_in_dma_address,               --                    Video_In_video_in_dma.address
			Video_In_video_in_dma_waitrequest              => video_in_video_in_dma_waitrequest,           --                                         .waitrequest
			Video_In_video_in_dma_write                    => video_in_video_in_dma_write,                 --                                         .write
			Video_In_video_in_dma_writedata                => video_in_video_in_dma_writedata,             --                                         .writedata
			Framebuffer_s1_address                         => mm_interconnect_0_framebuffer_s1_address,    --                           Framebuffer_s1.address
			Framebuffer_s1_write                           => mm_interconnect_0_framebuffer_s1_write,      --                                         .write
			Framebuffer_s1_readdata                        => mm_interconnect_0_framebuffer_s1_readdata,   --                                         .readdata
			Framebuffer_s1_writedata                       => mm_interconnect_0_framebuffer_s1_writedata,  --                                         .writedata
			Framebuffer_s1_chipselect                      => mm_interconnect_0_framebuffer_s1_chipselect, --                                         .chipselect
			Framebuffer_s1_clken                           => mm_interconnect_0_framebuffer_s1_clken       --                                         .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_50mhz_in_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of Raster_Laser_Projector
