-- Raster_Laser_Projector_X_Axis_Control.vhd

-- Generated using ACDS version 16.1 200

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Raster_Laser_Projector_X_Axis_Control is
	port (
		clk_in_clk             : in std_logic := '0'; --             clk_in.clk
		hsync_reference_in_clk : in std_logic := '0'; -- hsync_reference_in.clk
		reset_reset_n          : in std_logic := '0'; --              reset.reset_n
		reset_0_reset_n        : in std_logic := '0'  --            reset_0.reset_n
	);
end entity Raster_Laser_Projector_X_Axis_Control;

architecture rtl of Raster_Laser_Projector_X_Axis_Control is
begin

end architecture rtl; -- of Raster_Laser_Projector_X_Axis_Control
