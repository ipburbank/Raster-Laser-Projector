-- Raster_Laser_Projector_Video_In.vhd

-- Generated using ACDS version 16.1 200

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Raster_Laser_Projector_Video_In is
	port (
		clk_clk                                   : in  std_logic                     := '0';             --                         clk.clk
		reset_reset_n                             : in  std_logic                     := '0';             --                       reset.reset_n
		video_in_dma_address                      : out std_logic_vector(31 downto 0);                    --                video_in_dma.address
		video_in_dma_waitrequest                  : in  std_logic                     := '0';             --                            .waitrequest
		video_in_dma_write                        : out std_logic;                                        --                            .write
		video_in_dma_writedata                    : out std_logic_vector(7 downto 0);                     --                            .writedata
		video_in_external_interface_TD_CLK27      : in  std_logic                     := '0';             -- video_in_external_interface.TD_CLK27
		video_in_external_interface_TD_DATA       : in  std_logic_vector(7 downto 0)  := (others => '0'); --                            .TD_DATA
		video_in_external_interface_TD_HS         : in  std_logic                     := '0';             --                            .TD_HS
		video_in_external_interface_TD_VS         : in  std_logic                     := '0';             --                            .TD_VS
		video_in_external_interface_clk27_reset   : in  std_logic                     := '0';             --                            .clk27_reset
		video_in_external_interface_TD_RESET      : out std_logic;                                        --                            .TD_RESET
		video_in_external_interface_overflow_flag : out std_logic                                         --                            .overflow_flag
	);
end entity Raster_Laser_Projector_Video_In;

architecture rtl of Raster_Laser_Projector_Video_In is
	component Raster_Laser_Projector_Video_In_video_chroma_resampler_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component Raster_Laser_Projector_Video_In_video_chroma_resampler_0;

	component Raster_Laser_Projector_Video_In_video_clipper_0 is
		port (
			clk                      : in  std_logic                    := 'X';             -- clk
			reset                    : in  std_logic                    := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                    := 'X';             -- valid
			stream_in_ready          : out std_logic;                                       -- ready
			stream_out_ready         : in  std_logic                    := 'X';             -- ready
			stream_out_data          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                       -- startofpacket
			stream_out_endofpacket   : out std_logic;                                       -- endofpacket
			stream_out_valid         : out std_logic                                        -- valid
		);
	end component Raster_Laser_Projector_Video_In_video_clipper_0;

	component Raster_Laser_Projector_Video_In_video_csc is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component Raster_Laser_Projector_Video_In_video_csc;

	component Raster_Laser_Projector_Video_In_video_decoder_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0);                    -- data
			TD_CLK27                 : in  std_logic                     := 'X';             -- export
			TD_DATA                  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			TD_HS                    : in  std_logic                     := 'X';             -- export
			TD_VS                    : in  std_logic                     := 'X';             -- export
			clk27_reset              : in  std_logic                     := 'X';             -- export
			TD_RESET                 : out std_logic;                                        -- export
			overflow_flag            : out std_logic                                         -- export
		);
	end component Raster_Laser_Projector_Video_In_video_decoder_0;

	component Raster_Laser_Projector_Video_In_video_dma_controller_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(7 downto 0)                      -- writedata
		);
	end component Raster_Laser_Projector_Video_In_video_dma_controller_0;

	component Raster_Laser_Projector_Video_In_video_rgb_resampler_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component Raster_Laser_Projector_Video_In_video_rgb_resampler_0;

	component Raster_Laser_Projector_Video_In_video_scaler_0 is
		port (
			clk                      : in  std_logic                    := 'X';             -- clk
			reset                    : in  std_logic                    := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                    := 'X';             -- valid
			stream_in_ready          : out std_logic;                                       -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                    := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                       -- startofpacket
			stream_out_endofpacket   : out std_logic;                                       -- endofpacket
			stream_out_valid         : out std_logic;                                       -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_channel       : out std_logic                                        -- channel
		);
	end component Raster_Laser_Projector_Video_In_video_scaler_0;

	component Raster_Laser_Projector_Video_In_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                    := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                    := 'X';             -- reset
			in_0_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                    := 'X';             -- valid
			in_0_ready          : out std_logic;                                       -- ready
			in_0_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			in_0_channel        : in  std_logic                    := 'X';             -- channel
			out_0_data          : out std_logic_vector(7 downto 0);                    -- data
			out_0_valid         : out std_logic;                                       -- valid
			out_0_ready         : in  std_logic                    := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                       -- startofpacket
			out_0_endofpacket   : out std_logic                                        -- endofpacket
		);
	end component Raster_Laser_Projector_Video_In_avalon_st_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_clipper_0_avalon_clipper_source_valid           : std_logic;                     -- video_clipper_0:stream_out_valid -> video_scaler_0:stream_in_valid
	signal video_clipper_0_avalon_clipper_source_data            : std_logic_vector(7 downto 0);  -- video_clipper_0:stream_out_data -> video_scaler_0:stream_in_data
	signal video_clipper_0_avalon_clipper_source_ready           : std_logic;                     -- video_scaler_0:stream_in_ready -> video_clipper_0:stream_out_ready
	signal video_clipper_0_avalon_clipper_source_startofpacket   : std_logic;                     -- video_clipper_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	signal video_clipper_0_avalon_clipper_source_endofpacket     : std_logic;                     -- video_clipper_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	signal video_csc_avalon_csc_source_valid                     : std_logic;                     -- video_csc:stream_out_valid -> video_rgb_resampler_0:stream_in_valid
	signal video_csc_avalon_csc_source_data                      : std_logic_vector(23 downto 0); -- video_csc:stream_out_data -> video_rgb_resampler_0:stream_in_data
	signal video_csc_avalon_csc_source_ready                     : std_logic;                     -- video_rgb_resampler_0:stream_in_ready -> video_csc:stream_out_ready
	signal video_csc_avalon_csc_source_startofpacket             : std_logic;                     -- video_csc:stream_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	signal video_csc_avalon_csc_source_endofpacket               : std_logic;                     -- video_csc:stream_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	signal video_decoder_0_avalon_decoder_source_valid           : std_logic;                     -- video_decoder_0:stream_out_valid -> video_chroma_resampler_0:stream_in_valid
	signal video_decoder_0_avalon_decoder_source_data            : std_logic_vector(15 downto 0); -- video_decoder_0:stream_out_data -> video_chroma_resampler_0:stream_in_data
	signal video_decoder_0_avalon_decoder_source_ready           : std_logic;                     -- video_chroma_resampler_0:stream_in_ready -> video_decoder_0:stream_out_ready
	signal video_decoder_0_avalon_decoder_source_startofpacket   : std_logic;                     -- video_decoder_0:stream_out_startofpacket -> video_chroma_resampler_0:stream_in_startofpacket
	signal video_decoder_0_avalon_decoder_source_endofpacket     : std_logic;                     -- video_decoder_0:stream_out_endofpacket -> video_chroma_resampler_0:stream_in_endofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_valid         : std_logic;                     -- video_rgb_resampler_0:stream_out_valid -> video_clipper_0:stream_in_valid
	signal video_rgb_resampler_0_avalon_rgb_source_data          : std_logic_vector(7 downto 0);  -- video_rgb_resampler_0:stream_out_data -> video_clipper_0:stream_in_data
	signal video_rgb_resampler_0_avalon_rgb_source_ready         : std_logic;                     -- video_clipper_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	signal video_rgb_resampler_0_avalon_rgb_source_startofpacket : std_logic;                     -- video_rgb_resampler_0:stream_out_startofpacket -> video_clipper_0:stream_in_startofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_endofpacket   : std_logic;                     -- video_rgb_resampler_0:stream_out_endofpacket -> video_clipper_0:stream_in_endofpacket
	signal video_scaler_0_avalon_scaler_source_valid             : std_logic;                     -- video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	signal video_scaler_0_avalon_scaler_source_data              : std_logic_vector(7 downto 0);  -- video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	signal video_scaler_0_avalon_scaler_source_ready             : std_logic;                     -- avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	signal video_scaler_0_avalon_scaler_source_channel           : std_logic;                     -- video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	signal video_scaler_0_avalon_scaler_source_startofpacket     : std_logic;                     -- video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal video_scaler_0_avalon_scaler_source_endofpacket       : std_logic;                     -- video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                         : std_logic;                     -- avalon_st_adapter:out_0_valid -> video_dma_controller_0:stream_valid
	signal avalon_st_adapter_out_0_data                          : std_logic_vector(7 downto 0);  -- avalon_st_adapter:out_0_data -> video_dma_controller_0:stream_data
	signal avalon_st_adapter_out_0_ready                         : std_logic;                     -- video_dma_controller_0:stream_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                 : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> video_dma_controller_0:stream_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                   : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> video_dma_controller_0:stream_endofpacket
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, video_chroma_resampler_0:reset, video_clipper_0:reset, video_csc:reset, video_decoder_0:reset, video_dma_controller_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	signal reset_reset_n_ports_inv                               : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	video_chroma_resampler_0 : component Raster_Laser_Projector_Video_In_video_chroma_resampler_0
		port map (
			clk                      => clk_clk,                                             --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                      --                reset.reset
			stream_in_startofpacket  => video_decoder_0_avalon_decoder_source_startofpacket, --   avalon_chroma_sink.startofpacket
			stream_in_endofpacket    => video_decoder_0_avalon_decoder_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_decoder_0_avalon_decoder_source_valid,         --                     .valid
			stream_in_ready          => video_decoder_0_avalon_decoder_source_ready,         --                     .ready
			stream_in_data           => video_decoder_0_avalon_decoder_source_data,          --                     .data
			stream_out_ready         => open,                                                -- avalon_chroma_source.ready
			stream_out_startofpacket => open,                                                --                     .startofpacket
			stream_out_endofpacket   => open,                                                --                     .endofpacket
			stream_out_valid         => open,                                                --                     .valid
			stream_out_data          => open                                                 --                     .data
		);

	video_clipper_0 : component Raster_Laser_Projector_Video_In_video_clipper_0
		port map (
			clk                      => clk_clk,                                               --                   clk.clk
			reset                    => rst_controller_reset_out_reset,                        --                 reset.reset
			stream_in_data           => video_rgb_resampler_0_avalon_rgb_source_data,          --   avalon_clipper_sink.data
			stream_in_startofpacket  => video_rgb_resampler_0_avalon_rgb_source_startofpacket, --                      .startofpacket
			stream_in_endofpacket    => video_rgb_resampler_0_avalon_rgb_source_endofpacket,   --                      .endofpacket
			stream_in_valid          => video_rgb_resampler_0_avalon_rgb_source_valid,         --                      .valid
			stream_in_ready          => video_rgb_resampler_0_avalon_rgb_source_ready,         --                      .ready
			stream_out_ready         => video_clipper_0_avalon_clipper_source_ready,           -- avalon_clipper_source.ready
			stream_out_data          => video_clipper_0_avalon_clipper_source_data,            --                      .data
			stream_out_startofpacket => video_clipper_0_avalon_clipper_source_startofpacket,   --                      .startofpacket
			stream_out_endofpacket   => video_clipper_0_avalon_clipper_source_endofpacket,     --                      .endofpacket
			stream_out_valid         => video_clipper_0_avalon_clipper_source_valid            --                      .valid
		);

	video_csc : component Raster_Laser_Projector_Video_In_video_csc
		port map (
			clk                      => clk_clk,                                   --               clk.clk
			reset                    => rst_controller_reset_out_reset,            --             reset.reset
			stream_in_startofpacket  => open,                                      --   avalon_csc_sink.startofpacket
			stream_in_endofpacket    => open,                                      --                  .endofpacket
			stream_in_valid          => open,                                      --                  .valid
			stream_in_ready          => open,                                      --                  .ready
			stream_in_data           => open,                                      --                  .data
			stream_out_ready         => video_csc_avalon_csc_source_ready,         -- avalon_csc_source.ready
			stream_out_startofpacket => video_csc_avalon_csc_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_csc_avalon_csc_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_csc_avalon_csc_source_valid,         --                  .valid
			stream_out_data          => video_csc_avalon_csc_source_data           --                  .data
		);

	video_decoder_0 : component Raster_Laser_Projector_Video_In_video_decoder_0
		port map (
			clk                      => clk_clk,                                             --                   clk.clk
			reset                    => rst_controller_reset_out_reset,                      --                 reset.reset
			stream_out_ready         => video_decoder_0_avalon_decoder_source_ready,         -- avalon_decoder_source.ready
			stream_out_startofpacket => video_decoder_0_avalon_decoder_source_startofpacket, --                      .startofpacket
			stream_out_endofpacket   => video_decoder_0_avalon_decoder_source_endofpacket,   --                      .endofpacket
			stream_out_valid         => video_decoder_0_avalon_decoder_source_valid,         --                      .valid
			stream_out_data          => video_decoder_0_avalon_decoder_source_data,          --                      .data
			TD_CLK27                 => video_in_external_interface_TD_CLK27,                --    external_interface.export
			TD_DATA                  => video_in_external_interface_TD_DATA,                 --                      .export
			TD_HS                    => video_in_external_interface_TD_HS,                   --                      .export
			TD_VS                    => video_in_external_interface_TD_VS,                   --                      .export
			clk27_reset              => video_in_external_interface_clk27_reset,             --                      .export
			TD_RESET                 => video_in_external_interface_TD_RESET,                --                      .export
			overflow_flag            => video_in_external_interface_overflow_flag            --                      .export
		);

	video_dma_controller_0 : component Raster_Laser_Projector_Video_In_video_dma_controller_0
		port map (
			clk                  => clk_clk,                               --                      clk.clk
			reset                => rst_controller_reset_out_reset,        --                    reset.reset
			stream_data          => avalon_st_adapter_out_0_data,          --          avalon_dma_sink.data
			stream_startofpacket => avalon_st_adapter_out_0_startofpacket, --                         .startofpacket
			stream_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --                         .endofpacket
			stream_valid         => avalon_st_adapter_out_0_valid,         --                         .valid
			stream_ready         => avalon_st_adapter_out_0_ready,         --                         .ready
			slave_address        => open,                                  -- avalon_dma_control_slave.address
			slave_byteenable     => open,                                  --                         .byteenable
			slave_read           => open,                                  --                         .read
			slave_write          => open,                                  --                         .write
			slave_writedata      => open,                                  --                         .writedata
			slave_readdata       => open,                                  --                         .readdata
			master_address       => video_in_dma_address,                  --        avalon_dma_master.address
			master_waitrequest   => video_in_dma_waitrequest,              --                         .waitrequest
			master_write         => video_in_dma_write,                    --                         .write
			master_writedata     => video_in_dma_writedata                 --                         .writedata
		);

	video_rgb_resampler_0 : component Raster_Laser_Projector_Video_In_video_rgb_resampler_0
		port map (
			clk                      => clk_clk,                                               --               clk.clk
			reset                    => rst_controller_reset_out_reset,                        --             reset.reset
			stream_in_startofpacket  => video_csc_avalon_csc_source_startofpacket,             --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_csc_avalon_csc_source_endofpacket,               --                  .endofpacket
			stream_in_valid          => video_csc_avalon_csc_source_valid,                     --                  .valid
			stream_in_ready          => video_csc_avalon_csc_source_ready,                     --                  .ready
			stream_in_data           => video_csc_avalon_csc_source_data,                      --                  .data
			stream_out_ready         => video_rgb_resampler_0_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => video_rgb_resampler_0_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_rgb_resampler_0_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_rgb_resampler_0_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => video_rgb_resampler_0_avalon_rgb_source_data           --                  .data
		);

	video_scaler_0 : component Raster_Laser_Projector_Video_In_video_scaler_0
		port map (
			clk                      => clk_clk,                                             --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                      --                reset.reset
			stream_in_startofpacket  => video_clipper_0_avalon_clipper_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_clipper_0_avalon_clipper_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_clipper_0_avalon_clipper_source_valid,         --                     .valid
			stream_in_ready          => video_clipper_0_avalon_clipper_source_ready,         --                     .ready
			stream_in_data           => video_clipper_0_avalon_clipper_source_data,          --                     .data
			stream_out_ready         => video_scaler_0_avalon_scaler_source_ready,           -- avalon_scaler_source.ready
			stream_out_startofpacket => video_scaler_0_avalon_scaler_source_startofpacket,   --                     .startofpacket
			stream_out_endofpacket   => video_scaler_0_avalon_scaler_source_endofpacket,     --                     .endofpacket
			stream_out_valid         => video_scaler_0_avalon_scaler_source_valid,           --                     .valid
			stream_out_data          => video_scaler_0_avalon_scaler_source_data,            --                     .data
			stream_out_channel       => video_scaler_0_avalon_scaler_source_channel          --                     .channel
		);

	avalon_st_adapter : component Raster_Laser_Projector_Video_In_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 8,
			inChannelWidth  => 1,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                           -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,                    -- in_rst_0.reset
			in_0_data           => video_scaler_0_avalon_scaler_source_data,          --     in_0.data
			in_0_valid          => video_scaler_0_avalon_scaler_source_valid,         --         .valid
			in_0_ready          => video_scaler_0_avalon_scaler_source_ready,         --         .ready
			in_0_startofpacket  => video_scaler_0_avalon_scaler_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => video_scaler_0_avalon_scaler_source_endofpacket,   --         .endofpacket
			in_0_channel        => video_scaler_0_avalon_scaler_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_out_0_data,                      --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,                     --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,                     --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,             --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket                --         .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of Raster_Laser_Projector_Video_In
